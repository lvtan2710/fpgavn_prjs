////////////////////////////////////////////////////////////////////////////////
//
// FPGAVN.COM
//
// Filename     : a_fflopx.v
// Description  : This module is asynchronous flip-flop for a signal or a bus.
//
// Author       : fpgavn@fpgavn.com
// Created On   : Sat May 27 14:33:20 2017
// History (Date, Changed By)
//
////////////////////////////////////////////////////////////////////////////////

module a_fflopx.v
    (

     );

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations

////////////////////////////////////////////////////////////////////////////////
// Port declarations


////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation

endmodule 

////////////////////////////////////////////////////////////////////////////////
// 
// Company    : ROBERT BOSCH ENGINEERING VN
// Department : RBVH/EVH2
// Project    : 
// File       : a_fflopx.v
// Author     : Tan.LeVan@vn.bosch.com
// Created    : Wed Jul 15 19:18:36 2015
// Description: This module is asynchronous flip-flop for a signal or a bus.
// 
// History    : 
// 
////////////////////////////////////////////////////////////////////////////////

module a_fflopx
    (
     clk,
     rst_n,
     d,
     q
     );

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations
parameter           SIZE = 8;
parameter           RST_VAL = {SIZE{1'b0}};

////////////////////////////////////////////////////////////////////////////////
// Port declarations
input               clk;
input               rst_n;
input [SIZE-1:0]    d;
output [SIZE-1:0]   q;

////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation
reg [SIZE-1:0]      q;

always @(posedge clk or negedge rst_n)
    begin
    if (!rst_n) q <= RST_VAL;
    else        q <= d;
    end
    
endmodule 
