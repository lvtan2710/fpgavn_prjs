-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: alt_tdp_bram.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.0.0 Build 145 04/22/2015 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus II License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY alt_tdp_bram IS
  GENERIC (
    G_ADDR_A    : INTEGER := 10;
    G_WIDTH_A   : INTEGER := 16;
    G_DEPTH_A   : INTEGER := 1024;
    G_ADDR_B    : INTEGER := 10;
    G_WIDTH_B   : INTEGER := 16;
    G_DEPTH_B   : INTEGER := 1024;
    G_DEVICE    : STRING  := "zynq";
    G_COMMONCLK : INTEGER := 0;

    A_REG_EN_A  : STRING  := "CLOCK0";  -- CLOCK0, UNUSED
    A_REG_EN_B  : STRING  := "CLOCK1";  -- CLOCK0, CLOCK1, UNUSED
    A_WR_MODE   : STRING  := "NEW_DATA_NO_NBE_READ"; -- DONT_CARE, NEW_DATA_NO_NBE_READ
    A_MAXDEPTH  : INTEGER := 1024;
    A_BRAM_TYPE : STRING  := "AUTO"     -- AUTO, M512, M4K, M-RAM, MLAB, M9K, M144K, M10K, M20K, LC
                                        -- M512 blocks are not supported in true dual-port RAM mode
                                        -- MLAB blocks are not supported in simple dual-port RAM mode with mixed-width port feature, true dual-port RAM mode, and dual-port ROM mode 
    );
  PORT
	(
    address_a	: IN STD_LOGIC_VECTOR (G_ADDR_A-1 DOWNTO 0);
    address_b	: IN STD_LOGIC_VECTOR (G_ADDR_B-1 DOWNTO 0);
    data_a		: IN STD_LOGIC_VECTOR (G_WIDTH_A-1 DOWNTO 0);
    data_b		: IN STD_LOGIC_VECTOR (G_WIDTH_B-1 DOWNTO 0);
    inclock		: IN STD_LOGIC  := '1';
    outclock	: IN STD_LOGIC;
    wren_a		: IN STD_LOGIC  := '0';
    wren_b		: IN STD_LOGIC  := '0';
    q_a		    : OUT STD_LOGIC_VECTOR (G_WIDTH_A-1 DOWNTO 0);
    q_b		    : OUT STD_LOGIC_VECTOR (G_WIDTH_B-1 DOWNTO 0)
	);
END alt_tdp_bram;

ARCHITECTURE SYN OF alt_tdp_bram IS

  CONSTANT C_CLOCK0 : STRING := "CLOCK0";
  CONSTANT C_CLOCK1 : STRING := "CLOCK1";
  
  CONSTANT C_ADDRESS_REG_B : STRING := C_CLOCK1;-- := C_CLOCK0 WHEN (G_COMMONCLK = 1) ELSE C_CLOCK1;
  
  SIGNAL sub_wire0	: STD_LOGIC_VECTOR(G_WIDTH_A-1 DOWNTO 0);
  SIGNAL sub_wire1	: STD_LOGIC_VECTOR(G_WIDTH_B-1 DOWNTO 0);
  SIGNAL clock0     : STD_LOGIC;
  SIGNAL clock1     : STD_LOGIC;
    
BEGIN
	q_a    <= sub_wire0(G_WIDTH_A-1 DOWNTO 0);
	q_b    <= sub_wire1(G_WIDTH_B-1 DOWNTO 0);
    clock0 <= inclock;
    clock1 <= '1' WHEN (G_COMMONCLK = 1) ELSE outclock;
    
	altsyncram_component : altsyncram
	GENERIC MAP (
		address_reg_b           => C_ADDRESS_REG_B,
		clock_enable_input_a    => "BYPASS",
		clock_enable_input_b    => "BYPASS",
		clock_enable_output_a   => "BYPASS",
		clock_enable_output_b   => "BYPASS",
		indata_reg_b            => C_ADDRESS_REG_B,
		intended_device_family  => G_DEVICE,
		lpm_type                => "altsyncram",
        maximum_depth           => A_MAXDEPTH,
		numwords_a              => G_DEPTH_A,
		numwords_b              => G_DEPTH_B,
		operation_mode          => "BIDIR_DUAL_PORT",
		outdata_aclr_a          => "NONE",
		outdata_aclr_b          => "NONE",
		outdata_reg_a           => A_REG_EN_A,
		outdata_reg_b           => A_REG_EN_B,
		power_up_uninitialized  => "FALSE",
        ram_block_type          => A_BRAM_TYPE,
		read_during_write_mode_mixed_ports => "OLD_DATA",
		read_during_write_mode_port_a => A_WR_MODE,
		read_during_write_mode_port_b => A_WR_MODE,
		widthad_a               => G_ADDR_A,
		widthad_b               => G_ADDR_B,
		width_a                 => G_WIDTH_A,
		width_b                 => G_WIDTH_B,
		width_byteena_a         => 1,
		width_byteena_b         => 1,
		wrcontrol_wraddress_reg_b => C_ADDRESS_REG_B
	)
	PORT MAP (
		address_a   => address_a,
		address_b   => address_b,
		clock0      => clock0,
		clock1      => clock1,
		data_a      => data_a,
		data_b      => data_b,
		wren_a      => wren_a,
		wren_b      => wren_b,
		q_a         => sub_wire0,
		q_b         => sub_wire1
	);

END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_B NUMERIC "0"
-- Retrieval info: PRIVATE: CLRdata NUMERIC "0"
-- Retrieval info: PRIVATE: CLRq NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrren NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwren NUMERIC "0"
-- Retrieval info: PRIVATE: Clock NUMERIC "2"
-- Retrieval info: PRIVATE: Clock_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clock_B NUMERIC "0"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MEMSIZE NUMERIC "1024"
-- Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "3"
-- Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "1"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "3"
-- Retrieval info: PRIVATE: REGdata NUMERIC "1"
-- Retrieval info: PRIVATE: REGq NUMERIC "1"
-- Retrieval info: PRIVATE: REGrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: REGrren NUMERIC "0"
-- Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
-- Retrieval info: PRIVATE: REGwren NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
-- Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
-- Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
-- Retrieval info: PRIVATE: VarWidth NUMERIC "0"
-- Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "32"
-- Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "32"
-- Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "32"
-- Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "32"
-- Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: enable NUMERIC "0"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_B STRING "BYPASS"
-- Retrieval info: CONSTANT: INDATA_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "32"
-- Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "32"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "BIDIR_DUAL_PORT"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK1"
-- Retrieval info: CONSTANT: OUTDATA_REG_B STRING "CLOCK1"
-- Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_MIXED_PORTS STRING "OLD_DATA"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_A STRING "NEW_DATA_NO_NBE_READ"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_B STRING "NEW_DATA_NO_NBE_READ"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "5"
-- Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "5"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_B NUMERIC "1"
-- Retrieval info: CONSTANT: WRCONTROL_WRADDRESS_REG_B STRING "CLOCK0"
-- Retrieval info: USED_PORT: address_a 0 0 5 0 INPUT NODEFVAL "address_a[4..0]"
-- Retrieval info: USED_PORT: address_b 0 0 5 0 INPUT NODEFVAL "address_b[4..0]"
-- Retrieval info: USED_PORT: data_a 0 0 32 0 INPUT NODEFVAL "data_a[31..0]"
-- Retrieval info: USED_PORT: data_b 0 0 32 0 INPUT NODEFVAL "data_b[31..0]"
-- Retrieval info: USED_PORT: inclock 0 0 0 0 INPUT VCC "inclock"
-- Retrieval info: USED_PORT: outclock 0 0 0 0 INPUT NODEFVAL "outclock"
-- Retrieval info: USED_PORT: q_a 0 0 32 0 OUTPUT NODEFVAL "q_a[31..0]"
-- Retrieval info: USED_PORT: q_b 0 0 32 0 OUTPUT NODEFVAL "q_b[31..0]"
-- Retrieval info: USED_PORT: wren_a 0 0 0 0 INPUT GND "wren_a"
-- Retrieval info: USED_PORT: wren_b 0 0 0 0 INPUT GND "wren_b"
-- Retrieval info: CONNECT: @address_a 0 0 5 0 address_a 0 0 5 0
-- Retrieval info: CONNECT: @address_b 0 0 5 0 address_b 0 0 5 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 inclock 0 0 0 0
-- Retrieval info: CONNECT: @clock1 0 0 0 0 outclock 0 0 0 0
-- Retrieval info: CONNECT: @data_a 0 0 32 0 data_a 0 0 32 0
-- Retrieval info: CONNECT: @data_b 0 0 32 0 data_b 0 0 32 0
-- Retrieval info: CONNECT: @wren_a 0 0 0 0 wren_a 0 0 0 0
-- Retrieval info: CONNECT: @wren_b 0 0 0 0 wren_b 0 0 0 0
-- Retrieval info: CONNECT: q_a 0 0 32 0 @q_a 0 0 32 0
-- Retrieval info: CONNECT: q_b 0 0 32 0 @q_b 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_tdp_bram.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_tdp_bram.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_tdp_bram.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_tdp_bram.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_tdp_bram_inst.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_tdp_bram_syn.v TRUE
-- Retrieval info: LIB_FILE: altera_mf
