////////////////////////////////////////////////////////////////////////////////
//
// FPGAVN.COM
//
// Filename     : s_dff.v
// Description  : This module is a synchronous D-flipflop with low reset.
//
// Author       : fpgavn@fpgavn.com
// Created On   : Sat May 27 14:29:52 2017
// History (Date, Changed By)
//
////////////////////////////////////////////////////////////////////////////////

module s_dff
    (
     clk,
     rst_n,
     d,
     q
     );

////////////////////////////////////////////////////////////////////////////////
// Parameter declarations
parameter RST_VAL = 1'b0;

////////////////////////////////////////////////////////////////////////////////
// Port declarations
input     clk;
input     rst_n;
input     d;
output    q;

////////////////////////////////////////////////////////////////////////////////
// Local logic and instantiation
reg       q;
always @(posedge clk)
    begin
    if (!rst_n) q <= RST_VAL;
    else        q <= d;
    end
    
endmodule 
